`timescale 1ns / 1ps

module Solver_tb();


endmodule
